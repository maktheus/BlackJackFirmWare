module sevenSegmentes(
                    input wire [7:0] binario,
                    input wire clk,
                    output reg [7:0] seven_segments_signal_display
                    );

                    

endmodule