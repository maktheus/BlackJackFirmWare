module sevenSegmentes;

endmodule